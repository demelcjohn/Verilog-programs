module notgate(a, y);

input a;
output y;

not not1(y, a);

endmodule