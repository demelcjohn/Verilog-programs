module and2(x,y,out);

input x,y;
output out;

and and_gate(out,x,y);

endmodule
