module or2(x,y,out);

input x,y;
output out;

or or_gate(out,x,y);

endmodule
