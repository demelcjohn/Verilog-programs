module not1(x,out);
input x;
output out;
assign out = ~x;
endmodule
