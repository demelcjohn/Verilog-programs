module not2(x,out);

input x;
output out;

not not_gate(out,x);

endmodule
